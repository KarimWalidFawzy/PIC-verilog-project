module R_WCtrllgc(rdn,wrn,A0,CSn);
input rdn;


endmodule