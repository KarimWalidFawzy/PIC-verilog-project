module encode(
    input twotothen[0:7],
    output n[0:2]);


endmodule