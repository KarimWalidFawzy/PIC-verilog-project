module decode();
endmodule