module PRes();

endmodule