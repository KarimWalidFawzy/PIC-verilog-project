module CscdeCmprtr(CAS[0:2])
inout  CAS[0:2];

/*
1. 8259A outputs are master while the inputs are
slaves 
2.8259A (Master) sends the ID on CAS
3. Slave sends its routine 
*/
endmodule