module R_WCtrllgc(rdn,wrn,A0,CSn);
input rdn;
inout A0;
input wrn;
if(~(wrn|CSn))/** This detects pulses to see how to interact with 
CPU*/
if()


endmodule
